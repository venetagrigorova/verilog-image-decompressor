library verilog;
use verilog.vl_types.all;
entity tb_project_M1_v_unit is
end tb_project_M1_v_unit;
