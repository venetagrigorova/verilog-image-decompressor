library verilog;
use verilog.vl_types.all;
entity milestone1_v_unit is
end milestone1_v_unit;
