library verilog;
use verilog.vl_types.all;
entity milestone2_v_unit is
end milestone2_v_unit;
