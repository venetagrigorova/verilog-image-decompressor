library verilog;
use verilog.vl_types.all;
entity project_v_unit is
end project_v_unit;
